// ======== 7 Series ========
// AMD Spartan 7 Family
`define ID_7S6      32'h03622093
`define ID_7S15     32'h03620093
`define ID_7S25     32'h037C4093
`define ID_7S50     32'h0362F093
`define ID_7S75     32'h037C8093
`define ID_7S100    32'h037C7093

// AMD Artix 7 Family
`define ID_7A12T    32'h037C3093
`define ID_7A15T    32'h0362E093
`define ID_7A25T    32'h037C2093
`define ID_7A35T    32'h0362D093
`define ID_7A50T    32'h0362C093
`define ID_7A75T    32'h03632093
`define ID_7A100T   32'h03631093
`define ID_7A200T   32'h03636093

// AMD Kintex 7 Family
`define ID_7K70T    32'h03647093
`define ID_7K160T   32'h0364C093
`define ID_7K325T   32'h03651093
`define ID_7K355T   32'h03747093
`define ID_7K410T   32'h03656093
`define ID_7K420T   32'h03752093
`define ID_7K480T   32'h03751093

// AMD Virtex 7 Family
`define ID_7V585T   32'h03671093
`define ID_7V2000T  32'h036B3093
`define ID_7VX330T  32'h03667093
`define ID_7VX415T  32'h03682093
`define ID_7VX485T  32'h03687093
`define ID_7VX550T  32'h03692093
`define ID_7VX690T  32'h03691093
`define ID_7VX980T  32'h03696093
`define ID_7VX1140T 32'h036D5093
`define ID_7VH580T  32'h036D9093
`define ID_7VH870T  32'h036DB093

// ==== Ultrascale & Ultrascale+ ====
// Kintex UltraScale
`define ID_KU025    32'h03824093
`define ID_KU035    32'h03823093
`define ID_KU040    32'h03822093
`define ID_KU060    32'h03919093
`define ID_KU085    32'h0380F093
`define ID_KU095    32'h03844093
`define ID_KU115    32'h0390D093

// Virtex UltraScale
`define ID_VU065    32'h03939093
`define ID_VU080    32'h03843093
`define ID_VU095    32'h03842093
`define ID_VU125    32'h0392D093
`define ID_VU160    32'h03933093
`define ID_VU190    32'h03931093
`define ID_VU440    32'h0396D093

// Artix UltraScale+
`define ID_AU7P     32'h04AF6093
`define ID_AU10P    32'h04AC4093
`define ID_AU15P    32'h04AC2093
`define ID_AU20P    32'h04A65093
`define ID_AU25P    32'h04A64093

// Kintex UltraScale+
`define ID_KU3P     32'h04A63093
`define ID_KU5P     32'h04A62093
`define ID_KU9P     32'h0484A093
`define ID_KU11P    32'h04A4E093
`define ID_KU13P    32'h04A52093
`define ID_KU15P    32'h04A56093
`define ID_KU19P    32'h04ACF093

// Virtex UltraScale+
`define ID_VU3P     32'h04B39093
`define ID_VU5P     32'h04B2B093
`define ID_VU7P     32'h04B29093
`define ID_VU9P     32'h04B31093
`define ID_VU11P    32'h04B49093
`define ID_VU13P    32'h04B51093
`define ID_VU19P    32'h04BA1093
`define ID_VU23P    32'h04ACE093
`define ID_VU27P    32'h04B43093
`define ID_VU29P    32'h04B41093
`define ID_VU31P    32'h04B6B093
`define ID_VU33P    32'h04B69093
`define ID_VU35P    32'h04B71093
`define ID_VU37P    32'h04B79093
`define ID_VU45P    32'h04B73093
`define ID_VU47P    32'h04B7B093
`define ID_VU57P    32'h04B61093

